LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY IEEEtoBCD IS
	PORT(A:IN unsigned(63 downto 0);
		SBCD:OUT UNSIGNED(15 downto 0));
END ENTITY;

ARCHITECTURE comportamento OF IEEEtoBCD IS
	COMPONENT IEEEtoB is
		PORT (A:IN unsigned(62 DOWNTO 0);
			B: OUT unsigned(15 DOWNTO 0));
	END COMPONENT;
	COMPONENT BtoBCD IS
	PORT (A:IN UNSIGNED(15 DOWNTO 0);
		B: OUT UNSIGNED(15 DOWNTO 0));
	END COMPONENT;
	SIGNAL AUX1:unsigned(15 DOWNTO 0);
	BEGIN
	bc0:IEEEtoB PORT MAP(A(62 DOWNTO 0),AUX1);
	bc1:BtoBCD PORT MAP(AUX1,SBCD);



END ARCHITECTURE;

